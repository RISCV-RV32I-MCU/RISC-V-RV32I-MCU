module io_top
(
    input logic clk,
    input logic reset,
    // Bus Signals
    input logic bus_cs,
    input logic bus_wr,
    input logic bus_rd,
    input logic [31: 0] bus_addr,
    input logic [31: 0] bus_wr_data,
    output logic [31: 0] bus_rd_data,

    // UART
    input logic rx,
    output logic tx
    // SPI (optional)
            // input logic miso,
            // output logic sclk,
            // output logic mosi,
            // output logic ss_n
    // Matrix Multiplier
            //No IO
    // Cordic 
            //No IO
);

    // Register Declaration
    logic [15:0] mem_rd_array;
    logic [15:0] mem_wr_array;
    logic [15:0] cs_array;
    logic [4:0] reg_addr_array [16];
    logic [31:0] rd_data_array [16];
    logic [31:0] wr_data_array [16];

    // Instantiate I/O Controller
    io_controller ctrl_unit
    (
    .clk(clk),
    .reset(reset),
    .bus_cs(bus_cs),
    .bus_wr(bus_wr),
    .bus_rd(bus_rd),
    .bus_addr(bus_addr),
    .bus_wr_data(bus_wr_data),
    .bus_rd_data(bus_rd_data),
    // IO Slot Interface
    .slot_cs_array(cs_array),
    .slot_mem_rd_array(mem_rd_array),
    .slot_mem_wr_array(mem_wr_array),
    .slot_reg_addr_array(reg_addr_array),
    .slot_rd_data_array(rd_data_array),
    .slot_wr_data_array(wr_data_array)
    );

    // Slot 0: UART
    uart_top UART_MODULE
    (
    .clk(clk),
    .reset(reset),
    .cs(cs_array[0]),
    .read(mem_rd_array[0]),
    .write(mem_wr_array[0]),
    .addr(reg_addr_array[0]),
    .rd_data(rd_data_array[0]),
    .wr_data(wr_data_array[0]),

    .tx(tx),
    .rx(rx)
    );
    
    // Slot 1: Matrix Multiplier
    matrix_top MATRIX_MULTIPLIER_MODULE
    (
    .clk(clk),
    .reset(reset),
    .cs(cs_array[1]),
    .read(mem_rd_array[1]),
    .write(mem_wr_array[1]),
    .addr(reg_addr_array[1]),
    .rd_data(rd_data_array[1]),
    .wr_data(wr_data_array[1])
    );
    // Slot 2: Cordic Module
    cordic_top CORDIC_MODULE
    (
    .clk(clk),
    .reset(reset),
    .cs(cs_array[2]),
    .read(mem_rd_array[2]),
    .write(mem_wr_array[2]),
    .addr(reg_addr_array[2]),
    .rd_data(rd_data_array[2]),
    .wr_data(wr_data_array[2])
    );
    // Assign 0's to all unused slot rd_data signals
   generate
      genvar i;
       for (i=3; i<15; i=i+1) //Change as needed, this is assuming we used slots 0->2
        begin : gen_initialization_loop
            assign rd_data_array[i] = 32'h0;
        end
   endgenerate

endmodule
